package uart_env_pkg;
    import uvm_pkg::*;
    import uart_agent_pkg::*;
    import uart_ref_model_pkg::*;

    `include "uvm_macros.svh"
    `include "uart_scoreboard.sv"
    `include "uart_env.sv"
endpackage