package uart_ref_model_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import uart_agent_pkg::*;
    `include "uart_ref_model.sv"
endpackage