package uart_testlist_pkg;
    import uvm_pkg::*;
    import uart_env_pkg::*;
    import uart_seqlist_pkg::*;

    `include "uvm_macros.svh"
    `include "uart_basic_test.sv"
endpackage