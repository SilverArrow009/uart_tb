package uart_seqlist_pkg;
    import uvm_pkg::*;
    import uart_env_pkg::*;
    import uart_agent_pkg::*;
    
    `include "uvm_macros.svh"
    `include "uart_basic_sequence.sv"
endpackage